<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:demo="http://smartfrog.org/services/cdl/demo/">

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/cmp/components.cdl"/>

  <!--smartfrog extra classes-->

  <cdl:configuration>

    <!-- Echo something -->
    <demo:echo cdl:extends="cmp:Component">
      <cmp:CommandPath>
        org.smartfrog.services.cddlm.cdl.demo.EchoImpl</cmp:CommandPath>
      <demo:message sfi:type="trimmed"/>
      <demo:gui sfi:type="boolean">false</demo:gui>
    </demo:echo>


<!--    <demo:exec cdl:extends="cmp:Component">
      <cmp:CommandPath>
        org.smartfrog.services.cddlm.cdl.demo.JavaImpl</cmp:CommandPath>
    </demo:exec>-->


    <!--
    Run anything
    -->

    <demo:Run cdl:extends="cmp:Component">
      <cmp:CommandPath>
        org.smartfrog.services.os.runshell.RunShellImpl
      </cmp:CommandPath>

      <useExitCmd sfi:type="boolean">false</useExitCmd>
      <terminateOnFailure sfi:type="boolean">true</terminateOnFailure>
      <shouldTerminate sfi:type="boolean">true</shouldTerminate>
      <shellCmd sfi:type="trimmed"/>
      <exitCmd sfi:type="trimmed" sfi:optional="true"/>
      <workDir sfi:type="trimmed" sfi:optional="true"/>
      <logLevel sfi:type="integer">3</logLevel>
      <processID sfi:type="trimmed">demo:run</processID>
      <processName sfi:type="trimmed">demo:run</processName>
    </demo:Run>

    <!--Run Java -->
    <demo:Java cdl:extends="demo:Run">
      <classname sfi:type="trimmed"/>
      <jar sfi:type="trimmed"/>
      <maxMemory sfi:type="integer"/>
      <processID sfi:type="trimmed">demo:java</processID>
    </demo:Java>

    <demo:File cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.filesystem.FileImpl</cmp:CommandPath>
      <testOnDeploy sfi:type="boolean">false</testOnDeploy>
      <testOnLiveness sfi:type="boolean">true</testOnLiveness>
    </demo:File>

    <demo:Mkdir cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.filesystem.MkdirImpl</cmp:CommandPath>
      <dir sfi:type="trimmed"/>
      <parentDir sfi:type="trimmed" sfi:optional="true"/>
    </demo:Mkdir>


    <demo:TouchFile cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.filesystem.TouchFileImpl</cmp:CommandPath>
      <timestamp sfi:type="long">-1</timestamp>
    </demo:TouchFile>

    <demo:CopyFile cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.filesystem.CopyFileImpl</cmp:CommandPath>
      <source sfi:type="trimmed"/>
      <destination sfi:type="trimmed"/>
    </demo:CopyFile>

    <demo:DeployByCopy cdl:extends="demo:CopyFile">
      <cmp:CommandPath>org.smartfrog.services.filesystem.DeployByCopyImpl</cmp:CommandPath>
    </demo:DeployByCopy>

    <demo:TextFile cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.filesystem.TextFileImpl</cmp:CommandPath>
      <filename sfi:type="trimmed"/>
      <text sfi:type="string"/>
      <encoding sfi:type="UTF-8"/>
      <deleteOnExit sfi:type="boolean">false</deleteOnExit>
    </demo:TextFile>    
    
    <demo:Open cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.cddlm.cdl.demo.OpenImpl</cmp:CommandPath>
      <executable sfi:type="trimmed" sfi:optional="true" />
      <filename sfi:type="trimmed" sfi:optional="true"/>
    </demo:Open>
    
  </cdl:configuration>
</cdl:cdl>