<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:base="http://smartfrog.org/services/cdl/base/">


  <cdl:documentation>
    This set of components provides filesystem access
  </cdl:documentation>
  <!--smartfrog extra classes-->

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/base/components.cdl"/>

  <cdl:configuration>
  </cdl:configuration>
  <cdl:system>
    <composite cdl:extends="base:Compound"/>
  </cdl:system>
</cdl:cdl>

