<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
  xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
  xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
  xmlns:demo="http://smartfrog.org/services/cdl/demo/">

  <cdl:documentation>
    Echo something
  </cdl:documentation>
  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/demo/components.cdl"/>
  <cdl:configuration>
  </cdl:configuration>
  <cdl:system>
    <sfClass sfi:type="trimmed" cdl:ref="cmp:CommandPath"/>
    <cmp:CommandPath>org.smartfrog.services.cddlm.cdl.demo.EchoImpl</cmp:CommandPath>
    <demo:gui sfi:type="boolean">false</demo:gui>
    <demo:message sfi:type="trimmed">Test message</demo:message>
  </cdl:system>
</cdl:cdl>