<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:hosting="http://smartfrog.org/services/deployapi/components/hosting"
    >


  <cdl:documentation>
    This set of components represents some base classes of smartfrog, declared in CDL format
  </cdl:documentation>
  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/base/components.cdl"/>

  <cdl:configuration>

    <hosting:DeployapiCompound cdl:extends="base:Compound">
      <sfClass>org.smartfrog.services.deployapi.components.hosting.DeployapiCompoundImpl</sfClass>
    </hosting:DeployapiCompound>

  </cdl:configuration>
</cdl:cdl>