<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:demo="http://smartfrog.org/services/cdl/demo/">

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/cmp/components.cdl"/>

  <!--smartfrog extra classes-->

  <cdl:configuration>

    <!-- Echo something -->
    <demo:echo cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.cddlm.cdl.demo.EchoImpl</cmp:CommandPath>
      <demo:message sfi:type="trimmed"/>
      <demo:gui sfi:type="boolean">false</demo:gui>
    </demo:echo>


    <demo:exec cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.cddlm.cdl.demo.JavaImpl</cmp:CommandPath>
    </demo:exec>


    <demo:run cdl:extends="cmp:Component">
      <cmp:CommandPath>
        org.smartfrog.services.os.runshell.RunShellImpl
      </cmp:CommandPath>
      
      <useExitCmd sfi:type="boolean">false</useExitCmd>
      <terminateOnFailure sfi:type="boolean">true</terminateOnFailure>
      <shouldTerminate>true</shouldTerminate>
      <shellCmd sft:type="trimmed" />
      <exitCmd sft:type="trimmed"/>
      <logLevel sfi:type="int">3</logLevel>
      <processID sfi:type="trimmed">demo:run</processID>
    </demo:run>

  </cdl:configuration>
</cdl:cdl>