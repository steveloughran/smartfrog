<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="urn:cddlm/xml/0.1"
    xmlns:xs="http://www.w3.org/2001/XMLSchema"
    xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
    pathlanguage="http://w3c.org/"
    >
    <!--<import/>-->
    <cdl:types/>
    <cdl:configuration/>
    <cdl:system/>
</cdl:cdl>
