<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="urn:cddlm/xml/0.1"
    xmlns:xs="http://www.w3.org/2001/XMLSchema"
    xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
    >
    <cdl:system/>
    <cdl:configuration/>
    <cdl:types/>
</cdl:cdl>