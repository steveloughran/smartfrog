<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:base="http://smartfrog.org/services/cdl/base/">


  <cdl:documentation>
    Test for a lazy reference on a functional system.
    After deployment, app/user resolves to "lazy-value".
  </cdl:documentation>
  <!--smartfrog extra classes-->

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/base/components.cdl"/>

  <cdl:configuration>
    <toplevel>
      <value >lazy-value</value>
    </toplevel>
  </cdl:configuration>
  <cdl:system>
    <app>
      <user cdl:ref="value" cdl:lazy="true" cdl:refroot="toplevel"/>
    </app>
  </cdl:system>

</cdl:cdl>

