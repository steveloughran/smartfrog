<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:demo="http://smartfrog.org/services/cdl/demo/">

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/cmp/components.cdl"/>

  <!--smartfrog extra classes-->

  <cdl:configuration>

    <!-- Echo something -->
    <demo:echo cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.cddlm.cdl.demo.EchoImpl</cmp:CommandPath>
      <demo:message sfi:type="string"/>
      <demo:gui>false</demo:gui>
    </demo:echo>


    <demo:exec cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.cddlm.cdl.demo.JavaImpl</cmp:CommandPath>
    </demo:exec>


    <demo:java cdl:extends="cmp:Component">
      <cmp:CommandPath>
        org.smartfrog.services.cddlm.cdl.demo.CdlJavaImpl</cmp:CommandPath>
      <demo:classname />
    </demo:java>

  </cdl:configuration>
</cdl:cdl>