<?xml version="1.0"?>
<!-- this is not a valid CDL document -->
 <!-- the root element is of the wrong type -->
<cdl:types xmlns:cdl="http://gridforge.org/cddlm/xml/2004/07/30/"
    xmlns:xs="http://www.w3.org/2001/XMLSchema"
    xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
    >
</cdl:types>
