<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:base="http://smartfrog.org/services/cdl/base/">


  <cdl:documentation>
    This set of components provides filesystem access
  </cdl:documentation>
  <!--smartfrog extra classes-->

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/base/components.cdl"/>

  <cdl:configuration>


    <base:FileUsingComponent cdl:extends="base:Prim"/>


    <!--Declare the compound. sfSyncTerminate is trouble, as it is boolean not string-->
    <base:File cdl:extends="base:Prim">
      <sf:sfClass>org.smartfrog.services.filesystem.FileImpl</sf:sfClass>
    </base:File >

    <base:Mkdir cdl:extends="base:Prim">
      <sf:sfClass>org.smartfrog.services.filesystem.MkdirImpl</sf:sfClass>
    </base:Mkdir>


    <base:TempFile cdl:extends="base:FileUsingComponent">
      <sf:sfClass>org.smartfrog.services.filesystem.TempFile</sf:sfClass>
      <sf:encoding>UTF-8</sf:encoding>
      <sf:prefix>temp</sf:prefix>
      <sf:suffix>.tmp</sf:suffix>
<!--
      <sf:dir></sf:dir>
      <sf:text></sf:text>
-->
    </base:TempFile>


    <base:TouchFile cdl:extends="base:FileUsingComponent">
      <sf:sfClass>org.smartfrog.services.filesystem.TouchFileImpl</sf:sfClass>
    </base:TouchFile>

    <base:CopyFile cdl:extends="base:Compound">
      <sf:sfClass>org.smartfrog.services.filesystem.CopyFile</sf:sfClass>
<!--
      <sf:source />
      <sf:destination />
-->
    </base:CopyFile>

  </cdl:configuration>
</cdl:cdl>

