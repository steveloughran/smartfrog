<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:demo="http://smartfrog.org/services/cdl/demo/">


  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/demo/components.cdl"/>

  <cdl:configuration>
  </cdl:configuration>
  <cdl:system>
    <echo cdl:extends="demo:echo">
      <demo:message >
        Test message to antlai &amp; julgui
      </demo:message>
      <demo:gui>false</demo:gui>
    </echo>
  </cdl:system>
</cdl:cdl>

