<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://gridforge.org/cddlm/xml/2004/07/30/"
    xmlns:xs="http://www.w3.org/2001/XMLSchema"
    xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
  
    pathlanguage="http://w3c.org/"
    >
    <!--<import/>-->
    <cdl:types/>
    <cdl:configuration/>
    <cdl:system/>
</cdl:cdl>
