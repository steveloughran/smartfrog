<?xml version="1.0"?>
<!-- this is not a CDL document as it is not in the namespace -->
<cdl:cdl xmlns:cdl="urn:cddlm/xml/0.3"
    xmlns:xs="http://www.w3.org/2001/XMLSchema"
    xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
  xsi:schemaLocation="http://gridforge.org/cddlm/xml/2004/07/30/ cddlm.xsd"  
    >
    <!--<import/>-->
    <cdl:types>
    </cdl:types>
    <cdl:configuration xmlns="urn:other">


        <server cdl:name="server">
            <port>8080</port>
            <security>true</security>

            <webapps />
        </server>
        <server cdl:name="tomcat" cdl:extends="server">
            <basedir>
            </basedir>
        </server>

    </cdl:configuration>
    <cdl:system>
    </cdl:system>
</cdl:cdl>
