<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:demo="http://smartfrog.org/services/cdl/demo/"
    xmlns:jboss="http://smartfrog.org/services/cdl/demo/jboss">


  <cdl:documentation>
    This file defines JBoss and web components.
    It is not platform neutral, as it calls the shell/batch runtime to
    run different programs.
  </cdl:documentation>

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/demo/components.cdl"/>

  <cdl:configuration>

    <!--
         url extends OptionalString;
      //or
         //port of the page; default 80
         port extends OptionalInteger;
         //host of the page; default 127.0.0.1
         host extends OptionalString;
         //protocol, default http
         protocol extends OptionalString;
         //page
         page extends OptionalString;
         //query list of things that get turned into queries -without escaping.
         queries extends OptionalVector;

       //and any of

         //flag to set if you want any error text fetched from
         //the remote site. This is good for diagnostics.
         fetchErrorText extends OptionalBoolean;
         //response code below which the fetch is an error
         minimumResponseCode extends OptionalInteger;
         //error code above which an error has occurred,
         //default is 299.
         maximumResponseCode extends OptionalInteger;
         //flag to follow redirects
         followRedirects extends OptionalBoolean;
         //check frequency. This is the number of pings between checks
         //and so lets us probe less often than normal. default=1
         checkFrequency extends OptionalInteger;

         //flag to say that the check is on/off; useful during development
         enabled extends OptionalBoolean;

    -->
    <jboss:LivenessPage cdl:extends="cmp:Component">
      <sfClass>org.smartfrog.services.www.LivenessPageComponent</sfClass>
      <url sfi:type="trimmed" sfi:optional="true"/>
      <port sfi:type="integer" sfi:optional="true"/>
      <host sfi:type="trimmed" sfi:optional="true"/>
      <protocol sfi:type="trimmed" sfi:optional="true"/>
      <page sfi:type="trimmed" sfi:optional="true"/>
      <fetchErrorText sfi:type="boolean">true</fetchErrorText>
      <minimumResponseCode sfi:type="integer">200</minimumResponseCode>
      <maximumResponseCode sfi:type="integer">299</maximumResponseCode>
      <followRedirects sfi:type="boolean">true</followRedirects>
      <checkFrequency sfi:type="integer">1</checkFrequency>
    </jboss:LivenessPage>

    <jboss:JBoss cdl:extends="demo:Run">
      <homeDir sfi:type="trimmed"/>
      <deployDir sfi:type="trimmed"/>
      <processID>JBoss</processID>
      <!--bindings for the parent-->
      <workDir cdl:ref="homeDir"/>


    </jboss:JBoss>


    <jboss:JBossOnLinux cdl:extends="jboss:JBoss">
      <homeDir>/home/slo/jboss/</homeDir>
      <deployDir>/home/slo/jboss/server/default</deployDir>
      <shellCmd>/bin/bash /home/slo/jboss/bin/run.sh</shellCmd>
    </jboss:JBossOnLinux>

    <jboss:JBossOnDOS cdl:extends="jboss:JBoss">
      <homeDir>c:\Java\Apps\jboss-4.0\</homeDir>
      <deployDir>c:\Java\Apps\jboss-4.0\default</deployDir>
      <shellCmd>cmd.exe c:\Java\Apps\jboss-4.0\bin\run.bat</shellCmd>
    </jboss:JBossOnDOS>


    <jboss:System>

      <port>8080</port>
      <host>localhost</host>
      <application>diary</application>
      <source>c:\diary.war</source>

      <server cdl:extends="jboss:JBossOnDOS">
      </server>


      <jboss:demoWebApp cdl:extends="demo:DeployByCopy">
        <source cdl:ref="/source"/>
        <destination cdl:ref="/server/deployDir"/>
      </jboss:demoWebApp>


      <liveness cdl:extends="jboss:LivenessPage">
        <port cdl:ref="/port"/>
        <host cdl:ref="/host"/>
        <protocol>http</protocol>
        <page cdl:ref="/application"/>
      </liveness>


    </jboss:System>

  </cdl:configuration>


</cdl:cdl>