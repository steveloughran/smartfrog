<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="urn:cddlm/xml/0.1"
  xmlns:xs="http://www.w3.org/2001/XMLSchema"
  xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
  xsi:schemaLocation="urn:cddlm/xml/0.1 cddml.xsd">
  <!--<import/>-->
  <cdl:types/>
  <cdl:configuration>
    <cdl:component name="server">
      <port>8080</port>
      <security>true</security>
    </cdl:component>
    <cdl:component name="tomcat" extends="server">
      <basedir>
      </basedir>
    </cdl:component>

 </cdl:configuration>
  <cdl:system>
  </cdl:system>
</cdl:cdl>
